module restart